library verilog;
use verilog.vl_types.all;
entity combinational_circuit_vlg_check_tst is
    port(
        s1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end combinational_circuit_vlg_check_tst;
