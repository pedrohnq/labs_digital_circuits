library verilog;
use verilog.vl_types.all;
entity gates_vlg_check_tst is
    port(
        s1              : in     vl_logic;
        s2              : in     vl_logic;
        s3              : in     vl_logic;
        s4              : in     vl_logic;
        s5              : in     vl_logic;
        s6              : in     vl_logic;
        s7              : in     vl_logic;
        s8              : in     vl_logic;
        s9              : in     vl_logic;
        s10             : in     vl_logic;
        s11             : in     vl_logic;
        s12             : in     vl_logic;
        s13             : in     vl_logic;
        s14             : in     vl_logic;
        s15             : in     vl_logic;
        s16             : in     vl_logic;
        s17             : in     vl_logic;
        s18             : in     vl_logic;
        s19             : in     vl_logic;
        s20             : in     vl_logic;
        s21             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end gates_vlg_check_tst;
