library verilog;
use verilog.vl_types.all;
entity combinational_circuit_vlg_vec_tst is
end combinational_circuit_vlg_vec_tst;
