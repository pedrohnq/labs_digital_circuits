library verilog;
use verilog.vl_types.all;
entity gates is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        s1              : out    vl_logic;
        s2              : out    vl_logic;
        s3              : out    vl_logic;
        s4              : out    vl_logic;
        s5              : out    vl_logic;
        s6              : out    vl_logic;
        s7              : out    vl_logic;
        s8              : out    vl_logic;
        s9              : out    vl_logic;
        s10             : out    vl_logic;
        s11             : out    vl_logic;
        s12             : out    vl_logic;
        s13             : out    vl_logic;
        s14             : out    vl_logic;
        s15             : out    vl_logic;
        s16             : out    vl_logic;
        s17             : out    vl_logic;
        s18             : out    vl_logic;
        s19             : out    vl_logic;
        s20             : out    vl_logic;
        s21             : out    vl_logic
    );
end gates;
